vem bruno
